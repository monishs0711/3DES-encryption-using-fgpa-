module ip(input [1:64]M, output [1:32]L, output [33:64]R);
    wire [1:64] out;
    assign out[1] = M[58];
    assign out[2] = M[50];
    assign out[3] = M[42];
    assign out[4] = M[34];
    assign out[5] = M[26];
    assign out[6] = M[18];
    assign out[7] = M[10];
    assign out[8] = M[2];
    assign out[9] = M[60];
    assign out[10] = M[52];
    assign out[11] = M[44];
    assign out[12] = M[36];
    assign out[13] = M[28];
    assign out[14] = M[20];
    assign out[15] = M[12];
    assign out[16] = M[4];
    assign out[17] = M[62];
    assign out[18] = M[54];
    assign out[19] = M[46];
    assign out[20] = M[38];
    assign out[21] = M[30];
    assign out[22] = M[22];
    assign out[23] = M[14];
    assign out[24] = M[6];
    assign out[25] = M[64];
    assign out[26] = M[56];
    assign out[27] = M[48];
    assign out[28] = M[40];
    assign out[29] = M[32];
    assign out[30] = M[24];
    assign out[31] = M[16];
    assign out[32] = M[8];
    assign out[33] = M[57];
    assign out[34] = M[49];
    assign out[35] = M[41];
    assign out[36] = M[33];
    assign out[37] = M[25];
    assign out[38] = M[17];
    assign out[39] = M[9];
    assign out[40] = M[1];
    assign out[41] = M[59];
    assign out[42] = M[51];
    assign out[43] = M[43];
    assign out[44] = M[35];
    assign out[45] = M[27];
    assign out[46] = M[19];
    assign out[47] = M[11];
    assign out[48] = M[3];
    assign out[49] = M[61];
    assign out[50] = M[53];
    assign out[51] = M[45];
    assign out[52] = M[37];
    assign out[53] = M[29];
    assign out[54] = M[21];
    assign out[55] = M[13];
    assign out[56] = M[5];
    assign out[57] = M[63];
    assign out[58] = M[55];
    assign out[59] = M[47];
    assign out[60] = M[39];
    assign out[61] = M[31];
    assign out[62] = M[23];
    assign out[63] = M[15];
    assign out[64] = M[7];

    assign L = out[1:32];
    assign R = out[33:64];
endmodule