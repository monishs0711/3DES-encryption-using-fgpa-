module pc2 (input [1:28]c, [1:28]d ,output [1:48]subkey);
assign in={c,d};
assign subkey[1] = in[14];
assign subkey[2] = in[17];
assign subkey[3] = in[11];
assign subkey[4] = in[24];
assign subkey[5] = in[1];
assign subkey[6] = in[5];
assign subkey[7] = in[3];
assign subkey[8] = in[28];
assign subkey[9] = in[15];
assign subkey[10] = in[6];
assign subkey[11] = in[21];
assign subkey[12] = in[10];
assign subkey[13] = in[23];
assign subkey[14] = in[19];
assign subkey[15] = in[12];
assign subkey[16] = in[4];
assign subkey[17] = in[26];
assign subkey[18] = in[8];
assign subkey[19] = in[16];
assign subkey[20] = in[7];
assign subkey[21] = in[27];
assign subkey[22] = in[20];
assign subkey[23] = in[13];
assign subkey[24] = in[2];
assign subkey[25] = in[41];
assign subkey[26] = in[52];
assign subkey[27] = in[31];
assign subkey[28] = in[37];
assign subkey[29] = in[47];
assign subkey[30] = in[55];
assign subkey[31] = in[30];
assign subkey[32] = in[40];
assign subkey[33] = in[51];
assign subkey[34] = in[45];
assign subkey[35] = in[33];
assign subkey[36] = in[48];
assign subkey[37] = in[44];
assign subkey[38] = in[49];
assign subkey[39] = in[39];
assign subkey[40] = in[56];
assign subkey[41] = in[34];
assign subkey[42] = in[53];
assign subkey[43] = in[46];
assign subkey[44] = in[42];
assign subkey[45] = in[50];
assign subkey[46] = in[36];
assign subkey[47] = in[29];
assign subkey[48] = in[32];
endmodule